module MWCS(clk,reset,A,B,s,O);
input clk,reset,s;
input [31:0]A,B;
output [31:0]O;

wire [31:0]D[31:0];
wire [33:0]C0[9:0];
wire [33:0]S0[9:0];
wire [33:0]S0f;

wire [39:0]C1[5:0];
wire [39:0]S1[5:0];
wire [39:0]C1f[5:0];
wire [39:0]S1f[5:0];
wire [35:0]C16,C16f;
wire [35:0]S16,S16f;

wire [57:0]C2[3:0];
wire [57:0]S2[3:0];
wire [37:0]C24,C24f;
wire [37:0]S24;

wire [58:0]C3[1:0];
wire [58:0]S3[1:0];
wire [62:0]C32;
wire [62:0]S32;

wire [59:0]S40,C40;
wire [63:0]S41,C41;

wire [60:0]S5,C5;

wire [65:0]S6,C6;

wire [66:0]S70,C70;
wire [66:0]S71,C71;

wire [63:0]sum;

generate 
	genvar j,k;
	for(j=0; j<32; j=j+1) begin : AND_ROW
		for(k=0; k<32; k=k+1) begin : AND_Col
			and a0(D[j][k],A[k],B[j]);
		end
	end
endgenerate 

CSA #(34) c0({2'b00,D[0]},{1'b0,D[1],1'b0},{D[2],2'b00},S0[0],C0[0]);
CSA #(34) c1({2'b00,D[3]},{1'b0,D[4],1'b0},{D[5],2'b00},S0[1],C0[1]);
CSA #(34) c2({2'b00,D[6]},{1'b0,D[7],1'b0},{D[8],2'b00},S0[2],C0[2]);
CSA #(34) c3({2'b00,D[9]},{1'b0,D[10],1'b0},{D[11],2'b00},S0[3],C0[3]);
CSA #(34) c4({2'b00,D[12]},{1'b0,D[13],1'b0},{D[14],2'b00},S0[4],C0[4]);
CSA #(34) c5({2'b00,D[15]},{1'b0,D[16],1'b0},{D[17],2'b00},S0[5],C0[5]);
CSA #(34) c6({2'b00,D[18]},{1'b0,D[19],1'b0},{D[20],2'b00},S0[6],C0[6]);
CSA #(34) c7({2'b00,D[21]},{1'b0,D[22],1'b0},{D[23],2'b00},S0[7],C0[7]);
CSA #(34) c8({2'b00,D[24]},{1'b0,D[25],1'b0},{D[26],2'b00},S0[8],C0[8]);
CSA #(34) c9({2'b00,D[27]},{1'b0,D[28],1'b0},{D[29],2'b00},S0[9],C0[9]);

CSA #(40) c10({6'b0,S0[0]},{3'b0,S0[1],3'b0},{S0[2],6'b0},S1[0],C1[0]);
CSA #(40) c11({6'b0,S0[3]},{3'b0,S0[4],3'b0},{S0[5],6'b0},S1[1],C1[1]);
CSA #(40) c12({6'b0,S0[6]},{3'b0,S0[7],3'b0},{S0[8],6'b0},S1[2],C1[2]);
CSA #(40) c13({6'b0,C0[0]},{3'b0,C0[1],3'b0},{C0[2],6'b0},S1[3],C1[3]);
CSA #(40) c14({6'b0,C0[3]},{3'b0,C0[4],3'b0},{C0[5],6'b0},S1[4],C1[4]);
CSA #(40) c15({6'b0,C0[6]},{3'b0,C0[7],3'b0},{C0[8],6'b0},S1[5],C1[5]);
CSA #(36) c16({2'b0,C0[9]},{1'b0,D[30],3'b0},{D[31],4'b0},S16,C16);

FF32 #(586) ff1(clk,rset,{S1[0],S1[1],C1[0],C1[1],S1[2],S1[3],C1[2],C1[3],S1[4],S1[5],C1[4],C1[5],S16,C16,S0[9]}
        ,{S1f[0],S1f[1],C1f[0],C1f[1],S1f[2],S1f[3],C1f[2],C1f[3],S1f[4],S1f[5],C1f[4],C1f[5],S16f,C16f,S0f});

CSA #(58) c17({18'b0,S1f[0]},{9'b0,S1f[1],9'b0},{S1f[2],18'b0},S2[0],C2[0]);
CSA #(58) c18({18'b0,S1f[3]},{9'b0,S1f[4],9'b0},{S1f[5],18'b0},S2[1],C2[1]);
CSA #(58) c19({18'b0,C1f[0]},{9'b0,C1f[1],9'b0},{C1f[2],18'b0},S2[2],C2[2]);
CSA #(58) c20({18'b0,C1f[3]},{9'b0,C1f[4],9'b0},{C1f[5],18'b0},S2[3],C2[3]);
CSA #(38) c21({4'b0,S0f},{1'b0,S16f,1'b0},{C16f,2'b0},S24,C24);

CSA #(59) c22({1'b0,S2[0]},{S2[1],1'b0},{S2[2],1'b0},S3[0],C3[0]);
CSA #(59) c23({1'b0,C2[0]},{C2[1],1'b0},{C2[2],1'b0},S3[1],C3[1]);
CSA #(63) c24({5'b0,S2[3]},{4'b0,C2[3],1'b0},{S24,25'b0},S32,C32);

CSA #(60) c25({1'b0,S3[0]},{S3[1],1'b0},{C3[0],1'b0},S40,C40);
CSA #(64) c26({1'b0,S32},{C32,1'b0},{C24,26'b0},S41,C41);

CSA #(61) c27({1'b0,S40},{C40,1'b0},{C3[1],2'b0},S5,C5);

CSA #(66) c28({4'b0,S5},{S41,2'b0},{3'b0,C5,1'b0},S6,C6);

CSA #(67) c29({1'b0,S6},{C41,3'b0},{C6,26'b0},S70,C70);

FF32 #(134) ff2(clk,rset,{S70,C70},{S71,C71});

assign sum = S71[63:0] + C71[63:0];
assign O = (s)? sum[63:32] : sum[31:0];

endmodule 